import Vector::*;

typedef Vector#(pd, UInt#(pixelWidth)) Pixel#(numeric type pd, numeric type pixelWidth);
