`define IMPORT_HOSTIF 
`define XILINX_SYS_CLK 
`define ConnectalVersion 18.12.1
`define NumberOfMasters 1
`define PinType Top_Pins
`define PinTypeInclude Top_Pins
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 8
`define DerivedClockPeriod 10.000000
`define CnocTop 
`define XsimHostInterface 
`define PhysAddrWidth 40
`define SIMULATION 
`define CONNECTAL_BITS_DEPENDENCES bsim
`define BOARD_bluesim 
